import lc3b_types::*;

module ex_block
(
   input clk,
	input stall;
);

	  


endmodule : ex_block
