import lc3b_types::*;

module victim_cache
(
	input clk,

	
);


endmodule : victim_cache