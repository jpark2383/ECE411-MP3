import lc3b_types::*;

module mp3
(
    input clk,

    /* Memory signals */
    input pmem_resp,
    input logic[127:0] pmem_rdata,
    output pmem_read,
    output pmem_write,
    output lc3b_word pmem_address,
    output logic[127:0] pmem_wdata
);

	  


endmodule : mp3
