import lc3b_types::*;

module mem_block
(
   input clk,
	input stall;
);

	  


endmodule : mem_block
