import lc3b_types::*;

module datapath
(
    input clk,
    input stall,

);

	  


endmodule : datapath
